module bcd7seg(
  input  [3:0] b,
  output [7:0] h
);

    MuxKey #(16, 4, 8) i0 (h, b, {
        4'b0000, 8'b00000011,
        4'b0001, 8'b10011111,
        4'b0010, 8'b00100101,
        4'b0011, 8'b00001101,
        4'b0100, 8'b10011001,
        4'b0101, 8'b01001001,
        4'b0110, 8'b01000001,
        4'b0111, 8'b00011111,
        4'b1000, 8'b00000001,
        4'b1001, 8'b00001001,
        4'b1010, 8'b00010001,
        4'b1011, 8'b11000001,
        4'b1100, 8'b01100010,
        4'b1101, 8'b10000101,
        4'b1110, 8'b01100001,
        4'b1111, 8'b01110001
    });


endmodule

